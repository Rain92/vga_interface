`timescale 1ns / 1ns

module clock_converter_mmcme
  #(parameter MULT_F = 30.0, DIV_F = 25.0, DIVCLK_DIVIDE = 1,  CLKIN_PERIOD = 30.0)

   (
     input         clk_in,
     output        clk_out
   );

  wire clkfbout_buf;
  wire clkfbout;
  wire clk_out_;

  /* verilator lint_off PINCONNECTEMPTY */
  MMCME2_ADV
    #(.BANDWIDTH            ("OPTIMIZED"),
      .CLKOUT4_CASCADE      ("FALSE"),
      .COMPENSATION         ("ZHOLD"),
      .STARTUP_WAIT         ("FALSE"),
      .DIVCLK_DIVIDE        (DIVCLK_DIVIDE),
      .CLKFBOUT_MULT_F      (MULT_F),
      .CLKFBOUT_PHASE       (0.000),
      .CLKFBOUT_USE_FINE_PS ("FALSE"),
      .CLKOUT0_DIVIDE_F     (DIV_F),
      .CLKOUT0_PHASE        (0.000),
      .CLKOUT0_DUTY_CYCLE   (0.500),
      .CLKOUT0_USE_FINE_PS  ("FALSE"),
      .CLKIN1_PERIOD        (CLKIN_PERIOD))
    mmcm_adv_inst
    // Output clocks
    (
      .CLKFBOUT            (clkfbout),
      .CLKFBOUTB           (),
      .CLKOUT0             (clk_out_),
      .CLKOUT0B            (),
      .CLKOUT1             (),
      .CLKOUT1B            (),
      .CLKOUT2             (),
      .CLKOUT2B            (),
      .CLKOUT3             (),
      .CLKOUT3B            (),
      .CLKOUT4             (),
      .CLKOUT5             (),
      .CLKOUT6             (),
      // Input clock control
      .CLKFBIN             (clkfbout_buf),
      .CLKIN1              (clk_in),
      .CLKIN2              (1'b0),
      // Tied to always select the primary input clock
      .CLKINSEL            (1'b1),
      // Ports for dynamic reconfiguration
      .DADDR               (7'h0),
      .DCLK                (1'b0),
      .DEN                 (1'b0),
      .DI                  (16'h0),
      .DO                  (),
      .DRDY                (),
      .DWE                 (1'b0),
      // Ports for dynamic phase shift
      .PSCLK               (1'b0),
      .PSEN                (1'b0),
      .PSINCDEC            (1'b0),
      .PSDONE              (),
      // Other control and status signals
      .LOCKED              (),
      .CLKINSTOPPED        (),
      .CLKFBSTOPPED        (),
      .PWRDWN              (1'b0),
      .RST                 (1'b0));

  BUFG clkf_buf
       (.O (clkfbout_buf),
        .I (clkfbout));

  BUFG clkout1_buf
       (.O   (clk_out),
        .I   (clk_out_));

endmodule
